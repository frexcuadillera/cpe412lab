library verilog;
use verilog.vl_types.all;
entity demux18_behavioural_tb is
end demux18_behavioural_tb;

library verilog;
use verilog.vl_types.all;
entity synccntr3_tb is
end synccntr3_tb;

library verilog;
use verilog.vl_types.all;
entity demux18_dataflow_tb is
end demux18_dataflow_tb;

library verilog;
use verilog.vl_types.all;
entity mux21_tb is
end mux21_tb;

library verilog;
use verilog.vl_types.all;
entity VendingMoore_t is
end VendingMoore_t;

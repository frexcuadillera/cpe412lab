library verilog;
use verilog.vl_types.all;
entity mux81dataflow_tb is
end mux81dataflow_tb;

library verilog;
use verilog.vl_types.all;
entity dec_to_bin_encoder_tb is
end dec_to_bin_encoder_tb;

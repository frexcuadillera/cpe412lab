library verilog;
use verilog.vl_types.all;
entity jkff_tb is
end jkff_tb;

library verilog;
use verilog.vl_types.all;
entity mux41structural_tb is
end mux41structural_tb;

library verilog;
use verilog.vl_types.all;
entity sample_tb is
end sample_tb;

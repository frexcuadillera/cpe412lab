library verilog;
use verilog.vl_types.all;
entity decimal_to_priority_encoder_tb is
end decimal_to_priority_encoder_tb;

library verilog;
use verilog.vl_types.all;
entity mux81structural_tb is
end mux81structural_tb;

library verilog;
use verilog.vl_types.all;
entity \fa_tst_\ is
end \fa_tst_\;

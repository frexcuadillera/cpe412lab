library verilog;
use verilog.vl_types.all;
entity gated_d_latch_tb is
end gated_d_latch_tb;

`timescale 1ps/1ps
module jkff_tb();
  reg j,k,clk,reset;
  wire q;
  
  always #10 clk = ~clk;
  
  initial clk = 0;
  
  initial begin
    reset = 0;
  end
  
  initial begin
    {j,k} = 2'b11;
    #100 {j,k} = 2'b10;
  end
  
  initial begin
    #200
    {j,k} = 2'b11;
    #310 {j,k} = 2'b10;
  end
  
  initial begin
    #400
    {j,k} = 2'b11;
    #500 {j,k} = 2'b01;
  end
  
  initial begin
    #600
    {j,k} = 2'b11;
    #710 {j,k} = 2'b01;
  end
  
  initial begin
    #800 {j,k} = 2'b00;
    #1000 $stop;
  end
      
    jkff MUT(j,k,clk,reset,q);
    
endmodule                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   
library verilog;
use verilog.vl_types.all;
entity asynccnt3_tb is
end asynccnt3_tb;

library verilog;
use verilog.vl_types.all;
entity VendingMoore_tb is
end VendingMoore_tb;

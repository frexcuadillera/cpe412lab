library verilog;
use verilog.vl_types.all;
entity circuit_test is
end circuit_test;

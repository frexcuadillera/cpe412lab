module circuit(in1,in2,in3,in4,out);
  input in1,in2,in3,in4;
  output out;
  
  assign out = in1^in2^in3^in4;
  
  
endmodule

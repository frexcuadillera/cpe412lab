library verilog;
use verilog.vl_types.all;
entity magcomp2_tb is
end magcomp2_tb;

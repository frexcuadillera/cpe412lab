library verilog;
use verilog.vl_types.all;
entity master_slave_d_flip_flop_tb is
end master_slave_d_flip_flop_tb;
